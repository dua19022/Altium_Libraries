* BEGIN MODEL LME49860
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.  
*/////////////////////////////////////////////////////////////////////
* Legal Notice:  
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice. 
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND" 
*////////////////////////////////////////////////////////////////////
* PINOUT ORDER +IN -IN V+ V- OUT
* PINOUT ORDER  3   2   8  4  1
.SUBCKT LME49860 3 2 8 4 1
* NOTE THAT MODEL IS FOR ONE SECTION ONLY (A SECTION) OF
* THE DUAL LME49860
* MODEL FEATURES INCLUDE OUTPUT SWING, OUTPUT CURRENT THRU
* THE SUPPLY RAILS, OUTPUT CURRENT LIMIT, OPEN LOOP GAIN
* AND PHASE WITH CLOAD EFFECTS, SLEW RATE, COMMON MODE
* REJECTION WITH FREQ EFFECTS, POWER SUPPLY REJECTION WITH
* FREQ EFFECTS, INPUT VOLTAGE NOISE WITH 1/F, INPUT CURRENT
* NOISE WITH 1/F, INPUT BIAS CURRENT, OUTPUT IMPEDANCE,
* INPUT COMMON MODE RANGE, INPUT CAPACITANCE, INPUT OFFSET
* VOLTAGE WITH TEMPERATURE EFFECTS, AND QUIESCENT CURRENT
* VERSUS VOLTAGE.
* MODEL INCLUDES INPUT AND OUTPUT PROTECTION DIODES.
Q26 9 10 11 QON
Q27 12 10 13 QOP
Q28 4 14 15 QOP
Q29 8 16 17 QON
I4 9 16 3E-3
I5 14 12 3E-3
R34 18 17 1
R35 15 18 1
C6 10 19 2.8P
R36 19 10 1E3
G1 10 19 20 19 -1E-3
G2 21 19 22 23 -0.5E-2
R37 19 21 1.5E9
C7 20 24 15.33E-12
R38 20 21 1.9E3
E1 25 19 20 19 1
D2 25 21 DD
R39 19 24 45
Q30 23 26 27 QIN
Q31 22 28 29 QIN
Q32 30 31 32 QCN
R40 12 32 3.65E3
R41 23 33 220
R42 22 33 220
V7 9 34 0.75
R45 35 27 1
R46 35 29 1
R47 1 18 10
D1 34 33 DD
D3 21 25 DD
D4 36 9 DD
D5 12 37 DD
V8 36 21 1.5
V9 21 37 1.5
E6 38 0 9 0 1
E7 39 0 12 0 1
E8 40 0 41 0 1
R48 38 42 10E6
R49 39 43 10E6
R50 40 44 40E6
R51 0 42 10
R52 0 43 10
R53 0 44 40
E11 45 46 44 0 0.65
R54 47 41 1E3
R55 41 48 1E3
C10 38 42 1E-12
C11 39 43 1E-12
C12 40 44 0.4E-12
E12 49 45 43 0 0.30
E13 50 49 42 0 -0.62
R60 49 50 1E9
R61 45 49 1E9
R62 46 45 1E9
E22 47 0 2 0 1
E23 48 0 50 0 1
E24 51 52 53 54 17.5E-3
I7 0 54 1E-4
D6 54 0 DVN
I8 0 53 1E-4
D7 53 0 DVN
R63 26 50 19
R64 51 28 19
E25 12 0 4 0 1
E26 9 0 8 0 1
I9 8 4 5.8E-3
R65 4 8 19.23E3
E27 19 12 9 12 0.5
C13 2 0 3E-12
C14 50 0 3E-12
C15 50 2 0.25E-12
V10 52 2 87E-6
R67 13 16 1
R68 14 11 1
I13 50 0 -3.7313E-6
I14 2 0 -3.7313E-6
I15 12 31 3.442E-6
V12 35 30 -0.5
D8 55 26 DD
D9 55 28 DD
V13 55 12 1.45
I16 0 56 1E-3
D10 56 0 DD
R104 0 56 1E9
V14 56 57 0.65
R105 0 57 1E9
R106 0 57 1E9
E28 46 3 57 0 1.133E-4
R107 3 46 1E9
D11 26 9 DD
D12 28 9 DD
D13 1 58 DD
D14 59 1 DD
R108 58 8 10
R109 4 59 10
.MODEL DVN D KF=1.6E-13
.MODEL DD D
.MODEL QCN NPN
.MODEL QIN NPN BF=45 KF=2E-17
.MODEL QON NPN BF=15 RC=55
.MODEL QOP PNP BF=15 RC=55
.ENDS
* END MODEL LME49860
